VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_spraid
  CLASS BLOCK ;
  FOREIGN wrapped_spraid ;
  ORIGIN 0.000 0.000 ;
  SIZE 387.570 BY 398.290 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 394.290 51.110 398.290 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 67.740 387.570 68.940 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.270 0.000 249.830 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.230 0.000 261.790 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.350 0.000 386.910 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.390 0.000 374.950 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.150 0.000 124.710 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.100 4.000 70.300 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 164.300 387.570 165.500 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 103.100 387.570 104.300 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.190 0.000 273.750 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 394.290 158.750 398.290 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.030 0.000 344.590 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 270.380 387.570 271.580 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 394.290 98.950 398.290 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.670 394.290 337.230 398.290 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.780 4.000 325.980 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.670 394.290 360.230 398.290 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.550 394.290 212.110 398.290 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.790 0.000 255.350 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.940 4.000 62.140 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.830 0.000 220.390 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 394.290 116.430 398.290 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 394.290 63.070 398.290 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 394.290 140.350 398.290 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.860 4.000 194.060 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.470 0.000 351.030 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.510 0.000 178.070 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 85.420 387.570 86.620 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 394.290 21.670 398.290 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 243.180 387.570 244.380 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 0.000 285.710 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.980 4.000 387.180 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.190 0.000 112.750 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 0.000 148.630 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 0.000 279.270 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.300 4.000 97.500 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.260 4.000 44.460 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 0.000 225.910 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.350 394.290 294.910 398.290 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.110 0.000 297.670 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.310 394.290 306.870 398.290 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 209.180 387.570 210.380 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 305.740 387.570 306.940 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 199.660 387.570 200.860 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.500 4.000 158.700 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.550 0.000 166.110 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.150 394.290 354.710 398.290 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.780 4.000 87.980 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.990 0.000 356.550 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.900 4.000 9.100 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 0.000 95.270 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 357.420 387.570 358.620 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.710 394.290 325.270 398.290 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 0.000 29.950 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 0.000 107.230 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 191.500 387.570 192.700 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.390 0.000 213.950 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.980 4.000 149.180 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.110 394.290 205.670 398.290 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.620 4.000 351.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 394.290 81.470 398.290 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.070 394.290 378.630 398.290 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.990 394.290 241.550 398.290 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 331.580 387.570 332.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 341.100 387.570 342.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.380 4.000 237.580 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.230 394.290 330.790 398.290 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 226.860 387.570 228.060 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.350 394.290 110.910 398.290 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 59.580 387.570 60.780 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.140 4.000 395.340 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 394.290 86.990 398.290 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 366.940 387.570 368.140 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 156.140 387.570 157.340 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.070 394.290 33.630 398.290 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.060 4.000 17.260 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.950 0.000 184.510 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.540 4.000 211.740 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.390 394.290 259.950 398.290 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.590 394.290 384.150 398.290 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.260 4.000 316.460 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 0.000 35.470 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.670 394.290 176.230 398.290 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 32.380 387.570 33.580 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.190 394.290 342.750 398.290 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.580 4.000 26.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.180 4.000 176.380 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 0.000 291.230 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.630 394.290 372.190 398.290 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.870 394.290 277.430 398.290 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 217.340 387.570 218.540 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.780 4.000 359.980 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.070 0.000 332.630 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 128.940 387.570 130.140 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.950 394.290 253.510 398.290 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.790 394.290 301.350 398.290 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 77.260 387.570 78.460 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.430 394.290 270.990 398.290 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.270 394.290 134.830 398.290 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.630 394.290 188.190 398.290 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.470 394.290 236.030 398.290 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.550 0.000 327.110 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.430 0.000 362.990 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 0.000 53.870 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.220 4.000 263.420 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.030 394.290 229.590 398.290 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 138.460 387.570 139.660 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 14.700 387.570 15.900 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 394.290 39.150 398.290 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 323.420 387.570 324.620 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 386.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 386.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 386.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 386.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 386.480 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.710 394.290 164.270 398.290 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 384.620 387.570 385.820 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.100 4.000 342.300 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 235.020 387.570 236.220 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 313.900 387.570 315.100 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.900 4.000 281.100 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.430 0.000 17.990 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.590 0.000 131.150 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 41.900 387.570 43.100 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.510 394.290 224.070 398.290 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 0.000 155.070 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 6.540 387.570 7.740 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.110 0.000 320.670 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 394.290 16.150 398.290 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.100 4.000 308.300 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 181.980 387.570 183.180 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.460 4.000 377.660 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.660 4.000 166.860 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.070 0.000 309.630 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 394.290 152.310 398.290 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.110 0.000 136.670 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.860 4.000 228.060 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.580 4.000 298.780 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.820 4.000 141.020 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.230 394.290 146.790 398.290 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 0.000 100.790 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 394.290 93.430 398.290 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.950 0.000 368.510 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.430 0.000 201.990 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 296.220 387.570 297.420 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.420 4.000 52.620 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 0.000 83.310 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 394.290 122.870 398.290 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.750 0.000 267.310 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.420 4.000 290.620 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.270 394.290 318.830 398.290 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.990 394.290 57.550 398.290 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 394.290 128.390 398.290 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.110 394.290 182.670 398.290 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.150 394.290 170.710 398.290 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.990 0.000 11.550 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.830 0.000 59.390 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.300 4.000 131.500 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.030 0.000 160.590 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 375.100 387.570 376.300 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 394.290 69.510 398.290 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.070 394.290 217.630 398.290 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 0.000 41.910 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 94.940 387.570 96.140 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 278.540 387.570 279.740 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.700 4.000 219.900 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 173.820 387.570 175.020 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 394.290 9.710 398.290 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.620 4.000 79.820 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 349.260 387.570 350.460 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 394.290 247.990 398.290 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 0.000 88.830 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 112.620 387.570 113.820 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 0.000 237.870 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.910 0.000 380.470 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.550 394.290 28.110 398.290 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 0.000 303.190 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 0.000 47.430 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 0.000 143.110 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 50.060 387.570 51.260 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 392.780 387.570 393.980 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.140 4.000 123.340 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.590 0.000 315.150 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.340 4.000 184.540 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 120.780 387.570 121.980 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 0.000 6.030 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 288.060 387.570 289.260 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.110 394.290 366.670 398.290 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.510 0.000 339.070 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.710 394.290 348.270 398.290 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.060 4.000 255.260 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.740 4.000 272.940 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.870 0.000 208.430 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.830 0.000 243.390 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.940 4.000 334.140 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 394.290 75.030 398.290 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 394.290 200.150 398.290 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.540 4.000 245.740 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.270 0.000 65.830 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 0.000 23.510 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.910 394.290 265.470 398.290 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 394.290 193.710 398.290 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.990 0.000 172.550 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.750 394.290 313.310 398.290 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 24.220 387.570 25.420 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.300 4.000 369.500 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 260.860 387.570 262.060 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 0.000 71.350 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.630 0.000 119.190 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 0.000 190.030 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 252.700 387.570 253.900 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.910 0.000 196.470 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.830 394.290 289.390 398.290 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.390 394.290 282.950 398.290 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 394.290 45.590 398.290 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.830 394.290 105.390 398.290 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.620 4.000 113.820 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.630 394.290 4.190 398.290 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.570 146.620 387.570 147.820 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 7.225 385.335 386.325 ;
      LAYER met1 ;
        RECT 2.830 7.180 385.395 390.620 ;
      LAYER met2 ;
        RECT 0.090 394.010 3.350 394.925 ;
        RECT 4.470 394.010 8.870 394.925 ;
        RECT 9.990 394.010 15.310 394.925 ;
        RECT 16.430 394.010 20.830 394.925 ;
        RECT 21.950 394.010 27.270 394.925 ;
        RECT 28.390 394.010 32.790 394.925 ;
        RECT 33.910 394.010 38.310 394.925 ;
        RECT 39.430 394.010 44.750 394.925 ;
        RECT 45.870 394.010 50.270 394.925 ;
        RECT 51.390 394.010 56.710 394.925 ;
        RECT 57.830 394.010 62.230 394.925 ;
        RECT 63.350 394.010 68.670 394.925 ;
        RECT 69.790 394.010 74.190 394.925 ;
        RECT 75.310 394.010 80.630 394.925 ;
        RECT 81.750 394.010 86.150 394.925 ;
        RECT 87.270 394.010 92.590 394.925 ;
        RECT 93.710 394.010 98.110 394.925 ;
        RECT 99.230 394.010 104.550 394.925 ;
        RECT 105.670 394.010 110.070 394.925 ;
        RECT 111.190 394.010 115.590 394.925 ;
        RECT 116.710 394.010 122.030 394.925 ;
        RECT 123.150 394.010 127.550 394.925 ;
        RECT 128.670 394.010 133.990 394.925 ;
        RECT 135.110 394.010 139.510 394.925 ;
        RECT 140.630 394.010 145.950 394.925 ;
        RECT 147.070 394.010 151.470 394.925 ;
        RECT 152.590 394.010 157.910 394.925 ;
        RECT 159.030 394.010 163.430 394.925 ;
        RECT 164.550 394.010 169.870 394.925 ;
        RECT 170.990 394.010 175.390 394.925 ;
        RECT 176.510 394.010 181.830 394.925 ;
        RECT 182.950 394.010 187.350 394.925 ;
        RECT 188.470 394.010 192.870 394.925 ;
        RECT 193.990 394.010 199.310 394.925 ;
        RECT 200.430 394.010 204.830 394.925 ;
        RECT 205.950 394.010 211.270 394.925 ;
        RECT 212.390 394.010 216.790 394.925 ;
        RECT 217.910 394.010 223.230 394.925 ;
        RECT 224.350 394.010 228.750 394.925 ;
        RECT 229.870 394.010 235.190 394.925 ;
        RECT 236.310 394.010 240.710 394.925 ;
        RECT 241.830 394.010 247.150 394.925 ;
        RECT 248.270 394.010 252.670 394.925 ;
        RECT 253.790 394.010 259.110 394.925 ;
        RECT 260.230 394.010 264.630 394.925 ;
        RECT 265.750 394.010 270.150 394.925 ;
        RECT 271.270 394.010 276.590 394.925 ;
        RECT 277.710 394.010 282.110 394.925 ;
        RECT 283.230 394.010 288.550 394.925 ;
        RECT 289.670 394.010 294.070 394.925 ;
        RECT 295.190 394.010 300.510 394.925 ;
        RECT 301.630 394.010 306.030 394.925 ;
        RECT 307.150 394.010 312.470 394.925 ;
        RECT 313.590 394.010 317.990 394.925 ;
        RECT 319.110 394.010 324.430 394.925 ;
        RECT 325.550 394.010 329.950 394.925 ;
        RECT 331.070 394.010 336.390 394.925 ;
        RECT 337.510 394.010 341.910 394.925 ;
        RECT 343.030 394.010 347.430 394.925 ;
        RECT 348.550 394.010 353.870 394.925 ;
        RECT 354.990 394.010 359.390 394.925 ;
        RECT 360.510 394.010 365.830 394.925 ;
        RECT 366.950 394.010 371.350 394.925 ;
        RECT 372.470 394.010 377.790 394.925 ;
        RECT 378.910 394.010 383.310 394.925 ;
        RECT 0.090 4.280 384.000 394.010 ;
        RECT 0.790 4.000 5.190 4.280 ;
        RECT 6.310 4.000 10.710 4.280 ;
        RECT 11.830 4.000 17.150 4.280 ;
        RECT 18.270 4.000 22.670 4.280 ;
        RECT 23.790 4.000 29.110 4.280 ;
        RECT 30.230 4.000 34.630 4.280 ;
        RECT 35.750 4.000 41.070 4.280 ;
        RECT 42.190 4.000 46.590 4.280 ;
        RECT 47.710 4.000 53.030 4.280 ;
        RECT 54.150 4.000 58.550 4.280 ;
        RECT 59.670 4.000 64.990 4.280 ;
        RECT 66.110 4.000 70.510 4.280 ;
        RECT 71.630 4.000 76.950 4.280 ;
        RECT 78.070 4.000 82.470 4.280 ;
        RECT 83.590 4.000 87.990 4.280 ;
        RECT 89.110 4.000 94.430 4.280 ;
        RECT 95.550 4.000 99.950 4.280 ;
        RECT 101.070 4.000 106.390 4.280 ;
        RECT 107.510 4.000 111.910 4.280 ;
        RECT 113.030 4.000 118.350 4.280 ;
        RECT 119.470 4.000 123.870 4.280 ;
        RECT 124.990 4.000 130.310 4.280 ;
        RECT 131.430 4.000 135.830 4.280 ;
        RECT 136.950 4.000 142.270 4.280 ;
        RECT 143.390 4.000 147.790 4.280 ;
        RECT 148.910 4.000 154.230 4.280 ;
        RECT 155.350 4.000 159.750 4.280 ;
        RECT 160.870 4.000 165.270 4.280 ;
        RECT 166.390 4.000 171.710 4.280 ;
        RECT 172.830 4.000 177.230 4.280 ;
        RECT 178.350 4.000 183.670 4.280 ;
        RECT 184.790 4.000 189.190 4.280 ;
        RECT 190.310 4.000 195.630 4.280 ;
        RECT 196.750 4.000 201.150 4.280 ;
        RECT 202.270 4.000 207.590 4.280 ;
        RECT 208.710 4.000 213.110 4.280 ;
        RECT 214.230 4.000 219.550 4.280 ;
        RECT 220.670 4.000 225.070 4.280 ;
        RECT 226.190 4.000 231.510 4.280 ;
        RECT 232.630 4.000 237.030 4.280 ;
        RECT 238.150 4.000 242.550 4.280 ;
        RECT 243.670 4.000 248.990 4.280 ;
        RECT 250.110 4.000 254.510 4.280 ;
        RECT 255.630 4.000 260.950 4.280 ;
        RECT 262.070 4.000 266.470 4.280 ;
        RECT 267.590 4.000 272.910 4.280 ;
        RECT 274.030 4.000 278.430 4.280 ;
        RECT 279.550 4.000 284.870 4.280 ;
        RECT 285.990 4.000 290.390 4.280 ;
        RECT 291.510 4.000 296.830 4.280 ;
        RECT 297.950 4.000 302.350 4.280 ;
        RECT 303.470 4.000 308.790 4.280 ;
        RECT 309.910 4.000 314.310 4.280 ;
        RECT 315.430 4.000 319.830 4.280 ;
        RECT 320.950 4.000 326.270 4.280 ;
        RECT 327.390 4.000 331.790 4.280 ;
        RECT 332.910 4.000 338.230 4.280 ;
        RECT 339.350 4.000 343.750 4.280 ;
        RECT 344.870 4.000 350.190 4.280 ;
        RECT 351.310 4.000 355.710 4.280 ;
        RECT 356.830 4.000 362.150 4.280 ;
        RECT 363.270 4.000 367.670 4.280 ;
        RECT 368.790 4.000 374.110 4.280 ;
        RECT 375.230 4.000 379.630 4.280 ;
        RECT 380.750 4.000 384.000 4.280 ;
      LAYER met3 ;
        RECT 4.400 394.380 383.570 394.905 ;
        RECT 4.400 393.740 383.170 394.380 ;
        RECT 0.065 392.380 383.170 393.740 ;
        RECT 0.065 387.580 383.570 392.380 ;
        RECT 4.400 386.220 383.570 387.580 ;
        RECT 4.400 385.580 383.170 386.220 ;
        RECT 0.065 384.220 383.170 385.580 ;
        RECT 0.065 378.060 383.570 384.220 ;
        RECT 4.400 376.700 383.570 378.060 ;
        RECT 4.400 376.060 383.170 376.700 ;
        RECT 0.065 374.700 383.170 376.060 ;
        RECT 0.065 369.900 383.570 374.700 ;
        RECT 4.400 368.540 383.570 369.900 ;
        RECT 4.400 367.900 383.170 368.540 ;
        RECT 0.065 366.540 383.170 367.900 ;
        RECT 0.065 360.380 383.570 366.540 ;
        RECT 4.400 359.020 383.570 360.380 ;
        RECT 4.400 358.380 383.170 359.020 ;
        RECT 0.065 357.020 383.170 358.380 ;
        RECT 0.065 352.220 383.570 357.020 ;
        RECT 4.400 350.860 383.570 352.220 ;
        RECT 4.400 350.220 383.170 350.860 ;
        RECT 0.065 348.860 383.170 350.220 ;
        RECT 0.065 342.700 383.570 348.860 ;
        RECT 4.400 340.700 383.170 342.700 ;
        RECT 0.065 334.540 383.570 340.700 ;
        RECT 4.400 333.180 383.570 334.540 ;
        RECT 4.400 332.540 383.170 333.180 ;
        RECT 0.065 331.180 383.170 332.540 ;
        RECT 0.065 326.380 383.570 331.180 ;
        RECT 4.400 325.020 383.570 326.380 ;
        RECT 4.400 324.380 383.170 325.020 ;
        RECT 0.065 323.020 383.170 324.380 ;
        RECT 0.065 316.860 383.570 323.020 ;
        RECT 4.400 315.500 383.570 316.860 ;
        RECT 4.400 314.860 383.170 315.500 ;
        RECT 0.065 313.500 383.170 314.860 ;
        RECT 0.065 308.700 383.570 313.500 ;
        RECT 4.400 307.340 383.570 308.700 ;
        RECT 4.400 306.700 383.170 307.340 ;
        RECT 0.065 305.340 383.170 306.700 ;
        RECT 0.065 299.180 383.570 305.340 ;
        RECT 4.400 297.820 383.570 299.180 ;
        RECT 4.400 297.180 383.170 297.820 ;
        RECT 0.065 295.820 383.170 297.180 ;
        RECT 0.065 291.020 383.570 295.820 ;
        RECT 4.400 289.660 383.570 291.020 ;
        RECT 4.400 289.020 383.170 289.660 ;
        RECT 0.065 287.660 383.170 289.020 ;
        RECT 0.065 281.500 383.570 287.660 ;
        RECT 4.400 280.140 383.570 281.500 ;
        RECT 4.400 279.500 383.170 280.140 ;
        RECT 0.065 278.140 383.170 279.500 ;
        RECT 0.065 273.340 383.570 278.140 ;
        RECT 4.400 271.980 383.570 273.340 ;
        RECT 4.400 271.340 383.170 271.980 ;
        RECT 0.065 269.980 383.170 271.340 ;
        RECT 0.065 263.820 383.570 269.980 ;
        RECT 4.400 262.460 383.570 263.820 ;
        RECT 4.400 261.820 383.170 262.460 ;
        RECT 0.065 260.460 383.170 261.820 ;
        RECT 0.065 255.660 383.570 260.460 ;
        RECT 4.400 254.300 383.570 255.660 ;
        RECT 4.400 253.660 383.170 254.300 ;
        RECT 0.065 252.300 383.170 253.660 ;
        RECT 0.065 246.140 383.570 252.300 ;
        RECT 4.400 244.780 383.570 246.140 ;
        RECT 4.400 244.140 383.170 244.780 ;
        RECT 0.065 242.780 383.170 244.140 ;
        RECT 0.065 237.980 383.570 242.780 ;
        RECT 4.400 236.620 383.570 237.980 ;
        RECT 4.400 235.980 383.170 236.620 ;
        RECT 0.065 234.620 383.170 235.980 ;
        RECT 0.065 228.460 383.570 234.620 ;
        RECT 4.400 226.460 383.170 228.460 ;
        RECT 0.065 220.300 383.570 226.460 ;
        RECT 4.400 218.940 383.570 220.300 ;
        RECT 4.400 218.300 383.170 218.940 ;
        RECT 0.065 216.940 383.170 218.300 ;
        RECT 0.065 212.140 383.570 216.940 ;
        RECT 4.400 210.780 383.570 212.140 ;
        RECT 4.400 210.140 383.170 210.780 ;
        RECT 0.065 208.780 383.170 210.140 ;
        RECT 0.065 202.620 383.570 208.780 ;
        RECT 4.400 201.260 383.570 202.620 ;
        RECT 4.400 200.620 383.170 201.260 ;
        RECT 0.065 199.260 383.170 200.620 ;
        RECT 0.065 194.460 383.570 199.260 ;
        RECT 4.400 193.100 383.570 194.460 ;
        RECT 4.400 192.460 383.170 193.100 ;
        RECT 0.065 191.100 383.170 192.460 ;
        RECT 0.065 184.940 383.570 191.100 ;
        RECT 4.400 183.580 383.570 184.940 ;
        RECT 4.400 182.940 383.170 183.580 ;
        RECT 0.065 181.580 383.170 182.940 ;
        RECT 0.065 176.780 383.570 181.580 ;
        RECT 4.400 175.420 383.570 176.780 ;
        RECT 4.400 174.780 383.170 175.420 ;
        RECT 0.065 173.420 383.170 174.780 ;
        RECT 0.065 167.260 383.570 173.420 ;
        RECT 4.400 165.900 383.570 167.260 ;
        RECT 4.400 165.260 383.170 165.900 ;
        RECT 0.065 163.900 383.170 165.260 ;
        RECT 0.065 159.100 383.570 163.900 ;
        RECT 4.400 157.740 383.570 159.100 ;
        RECT 4.400 157.100 383.170 157.740 ;
        RECT 0.065 155.740 383.170 157.100 ;
        RECT 0.065 149.580 383.570 155.740 ;
        RECT 4.400 148.220 383.570 149.580 ;
        RECT 4.400 147.580 383.170 148.220 ;
        RECT 0.065 146.220 383.170 147.580 ;
        RECT 0.065 141.420 383.570 146.220 ;
        RECT 4.400 140.060 383.570 141.420 ;
        RECT 4.400 139.420 383.170 140.060 ;
        RECT 0.065 138.060 383.170 139.420 ;
        RECT 0.065 131.900 383.570 138.060 ;
        RECT 4.400 130.540 383.570 131.900 ;
        RECT 4.400 129.900 383.170 130.540 ;
        RECT 0.065 128.540 383.170 129.900 ;
        RECT 0.065 123.740 383.570 128.540 ;
        RECT 4.400 122.380 383.570 123.740 ;
        RECT 4.400 121.740 383.170 122.380 ;
        RECT 0.065 120.380 383.170 121.740 ;
        RECT 0.065 114.220 383.570 120.380 ;
        RECT 4.400 112.220 383.170 114.220 ;
        RECT 0.065 106.060 383.570 112.220 ;
        RECT 4.400 104.700 383.570 106.060 ;
        RECT 4.400 104.060 383.170 104.700 ;
        RECT 0.065 102.700 383.170 104.060 ;
        RECT 0.065 97.900 383.570 102.700 ;
        RECT 4.400 96.540 383.570 97.900 ;
        RECT 4.400 95.900 383.170 96.540 ;
        RECT 0.065 94.540 383.170 95.900 ;
        RECT 0.065 88.380 383.570 94.540 ;
        RECT 4.400 87.020 383.570 88.380 ;
        RECT 4.400 86.380 383.170 87.020 ;
        RECT 0.065 85.020 383.170 86.380 ;
        RECT 0.065 80.220 383.570 85.020 ;
        RECT 4.400 78.860 383.570 80.220 ;
        RECT 4.400 78.220 383.170 78.860 ;
        RECT 0.065 76.860 383.170 78.220 ;
        RECT 0.065 70.700 383.570 76.860 ;
        RECT 4.400 69.340 383.570 70.700 ;
        RECT 4.400 68.700 383.170 69.340 ;
        RECT 0.065 67.340 383.170 68.700 ;
        RECT 0.065 62.540 383.570 67.340 ;
        RECT 4.400 61.180 383.570 62.540 ;
        RECT 4.400 60.540 383.170 61.180 ;
        RECT 0.065 59.180 383.170 60.540 ;
        RECT 0.065 53.020 383.570 59.180 ;
        RECT 4.400 51.660 383.570 53.020 ;
        RECT 4.400 51.020 383.170 51.660 ;
        RECT 0.065 49.660 383.170 51.020 ;
        RECT 0.065 44.860 383.570 49.660 ;
        RECT 4.400 43.500 383.570 44.860 ;
        RECT 4.400 42.860 383.170 43.500 ;
        RECT 0.065 41.500 383.170 42.860 ;
        RECT 0.065 35.340 383.570 41.500 ;
        RECT 4.400 33.980 383.570 35.340 ;
        RECT 4.400 33.340 383.170 33.980 ;
        RECT 0.065 31.980 383.170 33.340 ;
        RECT 0.065 27.180 383.570 31.980 ;
        RECT 4.400 25.820 383.570 27.180 ;
        RECT 4.400 25.180 383.170 25.820 ;
        RECT 0.065 23.820 383.170 25.180 ;
        RECT 0.065 17.660 383.570 23.820 ;
        RECT 4.400 16.300 383.570 17.660 ;
        RECT 4.400 15.660 383.170 16.300 ;
        RECT 0.065 14.300 383.170 15.660 ;
        RECT 0.065 9.500 383.570 14.300 ;
        RECT 4.400 8.140 383.570 9.500 ;
        RECT 4.400 7.500 383.170 8.140 ;
        RECT 0.065 6.975 383.170 7.500 ;
      LAYER met4 ;
        RECT 0.295 17.855 20.640 373.145 ;
        RECT 23.040 17.855 97.440 373.145 ;
        RECT 99.840 17.855 174.240 373.145 ;
        RECT 176.640 17.855 251.040 373.145 ;
        RECT 253.440 17.855 327.840 373.145 ;
        RECT 330.240 17.855 370.465 373.145 ;
  END
END wrapped_spraid
END LIBRARY

