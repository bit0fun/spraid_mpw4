VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_spraid
  CLASS BLOCK ;
  FOREIGN wrapped_spraid ;
  ORIGIN 0.000 0.000 ;
  SIZE 397.755 BY 408.475 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.390 404.475 52.950 408.475 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 69.100 397.755 70.300 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 0.000 256.270 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.670 0.000 268.230 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 0.000 79.630 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.550 0.000 396.110 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.590 0.000 384.150 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 0.000 128.390 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.460 4.000 71.660 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 168.380 397.755 169.580 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 105.820 397.755 107.020 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.630 0.000 280.190 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 404.475 162.430 408.475 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 0.000 353.790 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 275.820 397.755 277.020 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.150 404.475 101.710 408.475 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.950 404.475 345.510 408.475 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.940 4.000 334.140 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.790 404.475 370.350 408.475 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.070 404.475 217.630 408.475 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.230 0.000 261.790 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 0.000 225.910 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.550 404.475 120.110 408.475 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 404.475 64.910 408.475 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 404.475 144.950 408.475 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.750 0.000 359.310 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.110 0.000 182.670 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 86.780 397.755 87.980 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.030 404.475 22.590 408.475 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 249.980 397.755 251.180 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.590 0.000 292.150 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.500 4.000 396.700 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 0.000 115.510 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 0.000 152.310 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 0.000 286.630 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.660 4.000 98.860 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.620 4.000 45.820 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.870 0.000 231.430 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 404.475 303.190 408.475 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.470 0.000 305.030 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.590 404.475 315.150 408.475 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 213.260 397.755 214.460 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 312.540 397.755 313.740 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 203.740 397.755 204.940 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.580 4.000 162.780 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.150 0.000 170.710 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.350 404.475 363.910 408.475 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.500 4.000 90.700 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 0.000 365.750 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.900 4.000 9.100 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 0.000 97.110 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 366.940 397.755 368.140 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.990 404.475 333.550 408.475 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 0.000 30.870 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 0.000 109.990 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 195.580 397.755 196.780 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 0.000 219.470 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.060 4.000 153.260 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 404.475 211.190 408.475 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.780 4.000 359.980 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 404.475 83.310 408.475 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.190 404.475 388.750 408.475 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 404.475 247.990 408.475 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 339.740 397.755 340.940 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 347.900 397.755 349.100 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.820 4.000 243.020 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 404.475 339.990 408.475 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 230.940 397.755 232.140 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 404.475 113.670 408.475 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 59.580 397.755 60.780 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.020 4.000 406.220 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.190 404.475 89.750 408.475 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 375.100 397.755 376.300 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 158.860 397.755 160.060 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.460 4.000 207.660 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 404.475 34.550 408.475 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.420 4.000 18.620 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.550 0.000 189.110 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.620 4.000 215.820 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 404.475 266.390 408.475 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.710 404.475 394.270 408.475 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.420 4.000 324.620 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.830 0.000 36.390 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 404.475 180.830 408.475 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 33.740 397.755 34.940 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 404.475 351.950 408.475 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.580 4.000 26.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.260 4.000 180.460 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 0.000 298.590 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.750 404.475 382.310 408.475 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.230 404.475 284.790 408.475 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 222.780 397.755 223.980 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.300 4.000 369.500 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.350 0.000 340.910 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 131.660 397.755 132.860 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.390 404.475 259.950 408.475 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.150 404.475 308.710 408.475 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 78.620 397.755 79.820 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.100 4.000 36.300 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.790 404.475 278.350 408.475 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 404.475 138.510 408.475 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 404.475 193.710 408.475 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.910 404.475 242.470 408.475 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.830 0.000 335.390 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.180 4.000 108.380 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.630 0.000 372.190 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.230 0.000 54.790 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.020 4.000 270.220 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.470 404.475 236.030 408.475 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 141.180 397.755 142.380 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 14.700 397.755 15.900 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 404.475 40.990 408.475 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 330.220 397.755 331.420 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 397.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 397.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 397.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 397.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 397.360 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.310 404.475 168.870 408.475 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 394.140 397.755 395.340 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.620 4.000 351.820 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 240.460 397.755 241.660 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 322.060 397.755 323.260 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.700 4.000 287.900 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.430 0.000 17.990 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 0.000 133.910 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 41.900 397.755 43.100 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.030 404.475 229.590 408.475 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 0.000 158.750 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 6.540 397.755 7.740 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.390 0.000 328.950 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.590 404.475 16.150 408.475 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.900 4.000 315.100 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 186.060 397.755 187.260 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.980 4.000 387.180 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.740 4.000 170.940 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.430 0.000 316.990 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 404.475 156.910 408.475 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 0.000 140.350 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.660 4.000 234.860 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.740 4.000 306.940 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.540 4.000 143.740 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.910 404.475 150.470 408.475 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 0.000 103.550 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 404.475 96.190 408.475 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 0.000 377.710 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.950 0.000 207.510 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 303.020 397.755 304.220 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.780 4.000 53.980 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.590 0.000 85.150 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 404.475 126.550 408.475 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.110 0.000 274.670 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.220 4.000 297.420 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.550 404.475 327.110 408.475 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.830 404.475 59.390 408.475 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.510 404.475 132.070 408.475 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 404.475 187.270 408.475 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 404.475 175.310 408.475 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.910 0.000 12.470 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 0.000 61.230 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.380 4.000 135.580 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.710 0.000 164.270 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 384.620 397.755 385.820 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 404.475 71.350 408.475 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.510 404.475 224.070 408.475 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 0.000 42.830 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 96.300 397.755 97.500 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 285.340 397.755 286.540 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.140 4.000 225.340 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 177.900 397.755 179.100 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.070 404.475 10.630 408.475 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.980 4.000 81.180 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 357.420 397.755 358.620 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.870 404.475 254.430 408.475 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 0.000 91.590 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 113.980 397.755 115.180 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.830 0.000 243.390 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 0.000 389.670 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 404.475 29.030 408.475 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 0.000 310.550 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.790 0.000 48.350 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 0.000 145.870 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 51.420 397.755 52.620 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 402.300 397.755 403.500 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.860 4.000 126.060 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.870 0.000 323.430 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 123.500 397.755 124.700 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 0.000 6.030 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 294.860 397.755 296.060 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.310 404.475 375.870 408.475 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.790 0.000 347.350 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.910 404.475 357.470 408.475 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.540 4.000 279.740 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 0.000 213.030 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.270 0.000 249.830 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.100 4.000 342.300 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 404.475 77.790 408.475 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.110 404.475 205.670 408.475 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.340 4.000 252.540 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.190 0.000 66.750 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.870 0.000 24.430 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.270 404.475 272.830 408.475 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 404.475 199.230 408.475 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 0.000 177.150 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.030 404.475 321.590 408.475 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 24.220 397.755 25.420 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.820 4.000 379.020 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 267.660 397.755 268.860 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 0.000 73.190 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 0.000 121.950 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.070 0.000 194.630 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 258.140 397.755 259.340 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.510 0.000 201.070 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.190 404.475 296.750 408.475 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 404.475 291.230 408.475 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 404.475 47.430 408.475 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.590 404.475 108.150 408.475 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 0.000 237.870 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.630 404.475 4.190 408.475 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.755 150.700 397.755 151.900 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 393.615 397.205 ;
      LAYER met1 ;
        RECT 0.070 7.520 394.150 397.360 ;
      LAYER met2 ;
        RECT 0.100 404.195 3.350 405.805 ;
        RECT 4.470 404.195 9.790 405.805 ;
        RECT 10.910 404.195 15.310 405.805 ;
        RECT 16.430 404.195 21.750 405.805 ;
        RECT 22.870 404.195 28.190 405.805 ;
        RECT 29.310 404.195 33.710 405.805 ;
        RECT 34.830 404.195 40.150 405.805 ;
        RECT 41.270 404.195 46.590 405.805 ;
        RECT 47.710 404.195 52.110 405.805 ;
        RECT 53.230 404.195 58.550 405.805 ;
        RECT 59.670 404.195 64.070 405.805 ;
        RECT 65.190 404.195 70.510 405.805 ;
        RECT 71.630 404.195 76.950 405.805 ;
        RECT 78.070 404.195 82.470 405.805 ;
        RECT 83.590 404.195 88.910 405.805 ;
        RECT 90.030 404.195 95.350 405.805 ;
        RECT 96.470 404.195 100.870 405.805 ;
        RECT 101.990 404.195 107.310 405.805 ;
        RECT 108.430 404.195 112.830 405.805 ;
        RECT 113.950 404.195 119.270 405.805 ;
        RECT 120.390 404.195 125.710 405.805 ;
        RECT 126.830 404.195 131.230 405.805 ;
        RECT 132.350 404.195 137.670 405.805 ;
        RECT 138.790 404.195 144.110 405.805 ;
        RECT 145.230 404.195 149.630 405.805 ;
        RECT 150.750 404.195 156.070 405.805 ;
        RECT 157.190 404.195 161.590 405.805 ;
        RECT 162.710 404.195 168.030 405.805 ;
        RECT 169.150 404.195 174.470 405.805 ;
        RECT 175.590 404.195 179.990 405.805 ;
        RECT 181.110 404.195 186.430 405.805 ;
        RECT 187.550 404.195 192.870 405.805 ;
        RECT 193.990 404.195 198.390 405.805 ;
        RECT 199.510 404.195 204.830 405.805 ;
        RECT 205.950 404.195 210.350 405.805 ;
        RECT 211.470 404.195 216.790 405.805 ;
        RECT 217.910 404.195 223.230 405.805 ;
        RECT 224.350 404.195 228.750 405.805 ;
        RECT 229.870 404.195 235.190 405.805 ;
        RECT 236.310 404.195 241.630 405.805 ;
        RECT 242.750 404.195 247.150 405.805 ;
        RECT 248.270 404.195 253.590 405.805 ;
        RECT 254.710 404.195 259.110 405.805 ;
        RECT 260.230 404.195 265.550 405.805 ;
        RECT 266.670 404.195 271.990 405.805 ;
        RECT 273.110 404.195 277.510 405.805 ;
        RECT 278.630 404.195 283.950 405.805 ;
        RECT 285.070 404.195 290.390 405.805 ;
        RECT 291.510 404.195 295.910 405.805 ;
        RECT 297.030 404.195 302.350 405.805 ;
        RECT 303.470 404.195 307.870 405.805 ;
        RECT 308.990 404.195 314.310 405.805 ;
        RECT 315.430 404.195 320.750 405.805 ;
        RECT 321.870 404.195 326.270 405.805 ;
        RECT 327.390 404.195 332.710 405.805 ;
        RECT 333.830 404.195 339.150 405.805 ;
        RECT 340.270 404.195 344.670 405.805 ;
        RECT 345.790 404.195 351.110 405.805 ;
        RECT 352.230 404.195 356.630 405.805 ;
        RECT 357.750 404.195 363.070 405.805 ;
        RECT 364.190 404.195 369.510 405.805 ;
        RECT 370.630 404.195 375.030 405.805 ;
        RECT 376.150 404.195 381.470 405.805 ;
        RECT 382.590 404.195 387.910 405.805 ;
        RECT 389.030 404.195 393.430 405.805 ;
        RECT 0.100 4.280 394.120 404.195 ;
        RECT 0.790 4.000 5.190 4.280 ;
        RECT 6.310 4.000 11.630 4.280 ;
        RECT 12.750 4.000 17.150 4.280 ;
        RECT 18.270 4.000 23.590 4.280 ;
        RECT 24.710 4.000 30.030 4.280 ;
        RECT 31.150 4.000 35.550 4.280 ;
        RECT 36.670 4.000 41.990 4.280 ;
        RECT 43.110 4.000 47.510 4.280 ;
        RECT 48.630 4.000 53.950 4.280 ;
        RECT 55.070 4.000 60.390 4.280 ;
        RECT 61.510 4.000 65.910 4.280 ;
        RECT 67.030 4.000 72.350 4.280 ;
        RECT 73.470 4.000 78.790 4.280 ;
        RECT 79.910 4.000 84.310 4.280 ;
        RECT 85.430 4.000 90.750 4.280 ;
        RECT 91.870 4.000 96.270 4.280 ;
        RECT 97.390 4.000 102.710 4.280 ;
        RECT 103.830 4.000 109.150 4.280 ;
        RECT 110.270 4.000 114.670 4.280 ;
        RECT 115.790 4.000 121.110 4.280 ;
        RECT 122.230 4.000 127.550 4.280 ;
        RECT 128.670 4.000 133.070 4.280 ;
        RECT 134.190 4.000 139.510 4.280 ;
        RECT 140.630 4.000 145.030 4.280 ;
        RECT 146.150 4.000 151.470 4.280 ;
        RECT 152.590 4.000 157.910 4.280 ;
        RECT 159.030 4.000 163.430 4.280 ;
        RECT 164.550 4.000 169.870 4.280 ;
        RECT 170.990 4.000 176.310 4.280 ;
        RECT 177.430 4.000 181.830 4.280 ;
        RECT 182.950 4.000 188.270 4.280 ;
        RECT 189.390 4.000 193.790 4.280 ;
        RECT 194.910 4.000 200.230 4.280 ;
        RECT 201.350 4.000 206.670 4.280 ;
        RECT 207.790 4.000 212.190 4.280 ;
        RECT 213.310 4.000 218.630 4.280 ;
        RECT 219.750 4.000 225.070 4.280 ;
        RECT 226.190 4.000 230.590 4.280 ;
        RECT 231.710 4.000 237.030 4.280 ;
        RECT 238.150 4.000 242.550 4.280 ;
        RECT 243.670 4.000 248.990 4.280 ;
        RECT 250.110 4.000 255.430 4.280 ;
        RECT 256.550 4.000 260.950 4.280 ;
        RECT 262.070 4.000 267.390 4.280 ;
        RECT 268.510 4.000 273.830 4.280 ;
        RECT 274.950 4.000 279.350 4.280 ;
        RECT 280.470 4.000 285.790 4.280 ;
        RECT 286.910 4.000 291.310 4.280 ;
        RECT 292.430 4.000 297.750 4.280 ;
        RECT 298.870 4.000 304.190 4.280 ;
        RECT 305.310 4.000 309.710 4.280 ;
        RECT 310.830 4.000 316.150 4.280 ;
        RECT 317.270 4.000 322.590 4.280 ;
        RECT 323.710 4.000 328.110 4.280 ;
        RECT 329.230 4.000 334.550 4.280 ;
        RECT 335.670 4.000 340.070 4.280 ;
        RECT 341.190 4.000 346.510 4.280 ;
        RECT 347.630 4.000 352.950 4.280 ;
        RECT 354.070 4.000 358.470 4.280 ;
        RECT 359.590 4.000 364.910 4.280 ;
        RECT 366.030 4.000 371.350 4.280 ;
        RECT 372.470 4.000 376.870 4.280 ;
        RECT 377.990 4.000 383.310 4.280 ;
        RECT 384.430 4.000 388.830 4.280 ;
        RECT 389.950 4.000 394.120 4.280 ;
      LAYER met3 ;
        RECT 4.400 404.620 393.755 405.785 ;
        RECT 4.000 403.900 393.755 404.620 ;
        RECT 4.000 401.900 393.355 403.900 ;
        RECT 4.000 397.100 393.755 401.900 ;
        RECT 4.400 395.740 393.755 397.100 ;
        RECT 4.400 395.100 393.355 395.740 ;
        RECT 4.000 393.740 393.355 395.100 ;
        RECT 4.000 387.580 393.755 393.740 ;
        RECT 4.400 386.220 393.755 387.580 ;
        RECT 4.400 385.580 393.355 386.220 ;
        RECT 4.000 384.220 393.355 385.580 ;
        RECT 4.000 379.420 393.755 384.220 ;
        RECT 4.400 377.420 393.755 379.420 ;
        RECT 4.000 376.700 393.755 377.420 ;
        RECT 4.000 374.700 393.355 376.700 ;
        RECT 4.000 369.900 393.755 374.700 ;
        RECT 4.400 368.540 393.755 369.900 ;
        RECT 4.400 367.900 393.355 368.540 ;
        RECT 4.000 366.540 393.355 367.900 ;
        RECT 4.000 360.380 393.755 366.540 ;
        RECT 4.400 359.020 393.755 360.380 ;
        RECT 4.400 358.380 393.355 359.020 ;
        RECT 4.000 357.020 393.355 358.380 ;
        RECT 4.000 352.220 393.755 357.020 ;
        RECT 4.400 350.220 393.755 352.220 ;
        RECT 4.000 349.500 393.755 350.220 ;
        RECT 4.000 347.500 393.355 349.500 ;
        RECT 4.000 342.700 393.755 347.500 ;
        RECT 4.400 341.340 393.755 342.700 ;
        RECT 4.400 340.700 393.355 341.340 ;
        RECT 4.000 339.340 393.355 340.700 ;
        RECT 4.000 334.540 393.755 339.340 ;
        RECT 4.400 332.540 393.755 334.540 ;
        RECT 4.000 331.820 393.755 332.540 ;
        RECT 4.000 329.820 393.355 331.820 ;
        RECT 4.000 325.020 393.755 329.820 ;
        RECT 4.400 323.660 393.755 325.020 ;
        RECT 4.400 323.020 393.355 323.660 ;
        RECT 4.000 321.660 393.355 323.020 ;
        RECT 4.000 315.500 393.755 321.660 ;
        RECT 4.400 314.140 393.755 315.500 ;
        RECT 4.400 313.500 393.355 314.140 ;
        RECT 4.000 312.140 393.355 313.500 ;
        RECT 4.000 307.340 393.755 312.140 ;
        RECT 4.400 305.340 393.755 307.340 ;
        RECT 4.000 304.620 393.755 305.340 ;
        RECT 4.000 302.620 393.355 304.620 ;
        RECT 4.000 297.820 393.755 302.620 ;
        RECT 4.400 296.460 393.755 297.820 ;
        RECT 4.400 295.820 393.355 296.460 ;
        RECT 4.000 294.460 393.355 295.820 ;
        RECT 4.000 288.300 393.755 294.460 ;
        RECT 4.400 286.940 393.755 288.300 ;
        RECT 4.400 286.300 393.355 286.940 ;
        RECT 4.000 284.940 393.355 286.300 ;
        RECT 4.000 280.140 393.755 284.940 ;
        RECT 4.400 278.140 393.755 280.140 ;
        RECT 4.000 277.420 393.755 278.140 ;
        RECT 4.000 275.420 393.355 277.420 ;
        RECT 4.000 270.620 393.755 275.420 ;
        RECT 4.400 269.260 393.755 270.620 ;
        RECT 4.400 268.620 393.355 269.260 ;
        RECT 4.000 267.260 393.355 268.620 ;
        RECT 4.000 262.460 393.755 267.260 ;
        RECT 4.400 260.460 393.755 262.460 ;
        RECT 4.000 259.740 393.755 260.460 ;
        RECT 4.000 257.740 393.355 259.740 ;
        RECT 4.000 252.940 393.755 257.740 ;
        RECT 4.400 251.580 393.755 252.940 ;
        RECT 4.400 250.940 393.355 251.580 ;
        RECT 4.000 249.580 393.355 250.940 ;
        RECT 4.000 243.420 393.755 249.580 ;
        RECT 4.400 242.060 393.755 243.420 ;
        RECT 4.400 241.420 393.355 242.060 ;
        RECT 4.000 240.060 393.355 241.420 ;
        RECT 4.000 235.260 393.755 240.060 ;
        RECT 4.400 233.260 393.755 235.260 ;
        RECT 4.000 232.540 393.755 233.260 ;
        RECT 4.000 230.540 393.355 232.540 ;
        RECT 4.000 225.740 393.755 230.540 ;
        RECT 4.400 224.380 393.755 225.740 ;
        RECT 4.400 223.740 393.355 224.380 ;
        RECT 4.000 222.380 393.355 223.740 ;
        RECT 4.000 216.220 393.755 222.380 ;
        RECT 4.400 214.860 393.755 216.220 ;
        RECT 4.400 214.220 393.355 214.860 ;
        RECT 4.000 212.860 393.355 214.220 ;
        RECT 4.000 208.060 393.755 212.860 ;
        RECT 4.400 206.060 393.755 208.060 ;
        RECT 4.000 205.340 393.755 206.060 ;
        RECT 4.000 203.340 393.355 205.340 ;
        RECT 4.000 198.540 393.755 203.340 ;
        RECT 4.400 197.180 393.755 198.540 ;
        RECT 4.400 196.540 393.355 197.180 ;
        RECT 4.000 195.180 393.355 196.540 ;
        RECT 4.000 190.380 393.755 195.180 ;
        RECT 4.400 188.380 393.755 190.380 ;
        RECT 4.000 187.660 393.755 188.380 ;
        RECT 4.000 185.660 393.355 187.660 ;
        RECT 4.000 180.860 393.755 185.660 ;
        RECT 4.400 179.500 393.755 180.860 ;
        RECT 4.400 178.860 393.355 179.500 ;
        RECT 4.000 177.500 393.355 178.860 ;
        RECT 4.000 171.340 393.755 177.500 ;
        RECT 4.400 169.980 393.755 171.340 ;
        RECT 4.400 169.340 393.355 169.980 ;
        RECT 4.000 167.980 393.355 169.340 ;
        RECT 4.000 163.180 393.755 167.980 ;
        RECT 4.400 161.180 393.755 163.180 ;
        RECT 4.000 160.460 393.755 161.180 ;
        RECT 4.000 158.460 393.355 160.460 ;
        RECT 4.000 153.660 393.755 158.460 ;
        RECT 4.400 152.300 393.755 153.660 ;
        RECT 4.400 151.660 393.355 152.300 ;
        RECT 4.000 150.300 393.355 151.660 ;
        RECT 4.000 144.140 393.755 150.300 ;
        RECT 4.400 142.780 393.755 144.140 ;
        RECT 4.400 142.140 393.355 142.780 ;
        RECT 4.000 140.780 393.355 142.140 ;
        RECT 4.000 135.980 393.755 140.780 ;
        RECT 4.400 133.980 393.755 135.980 ;
        RECT 4.000 133.260 393.755 133.980 ;
        RECT 4.000 131.260 393.355 133.260 ;
        RECT 4.000 126.460 393.755 131.260 ;
        RECT 4.400 125.100 393.755 126.460 ;
        RECT 4.400 124.460 393.355 125.100 ;
        RECT 4.000 123.100 393.355 124.460 ;
        RECT 4.000 118.300 393.755 123.100 ;
        RECT 4.400 116.300 393.755 118.300 ;
        RECT 4.000 115.580 393.755 116.300 ;
        RECT 4.000 113.580 393.355 115.580 ;
        RECT 4.000 108.780 393.755 113.580 ;
        RECT 4.400 107.420 393.755 108.780 ;
        RECT 4.400 106.780 393.355 107.420 ;
        RECT 4.000 105.420 393.355 106.780 ;
        RECT 4.000 99.260 393.755 105.420 ;
        RECT 4.400 97.900 393.755 99.260 ;
        RECT 4.400 97.260 393.355 97.900 ;
        RECT 4.000 95.900 393.355 97.260 ;
        RECT 4.000 91.100 393.755 95.900 ;
        RECT 4.400 89.100 393.755 91.100 ;
        RECT 4.000 88.380 393.755 89.100 ;
        RECT 4.000 86.380 393.355 88.380 ;
        RECT 4.000 81.580 393.755 86.380 ;
        RECT 4.400 80.220 393.755 81.580 ;
        RECT 4.400 79.580 393.355 80.220 ;
        RECT 4.000 78.220 393.355 79.580 ;
        RECT 4.000 72.060 393.755 78.220 ;
        RECT 4.400 70.700 393.755 72.060 ;
        RECT 4.400 70.060 393.355 70.700 ;
        RECT 4.000 68.700 393.355 70.060 ;
        RECT 4.000 63.900 393.755 68.700 ;
        RECT 4.400 61.900 393.755 63.900 ;
        RECT 4.000 61.180 393.755 61.900 ;
        RECT 4.000 59.180 393.355 61.180 ;
        RECT 4.000 54.380 393.755 59.180 ;
        RECT 4.400 53.020 393.755 54.380 ;
        RECT 4.400 52.380 393.355 53.020 ;
        RECT 4.000 51.020 393.355 52.380 ;
        RECT 4.000 46.220 393.755 51.020 ;
        RECT 4.400 44.220 393.755 46.220 ;
        RECT 4.000 43.500 393.755 44.220 ;
        RECT 4.000 41.500 393.355 43.500 ;
        RECT 4.000 36.700 393.755 41.500 ;
        RECT 4.400 35.340 393.755 36.700 ;
        RECT 4.400 34.700 393.355 35.340 ;
        RECT 4.000 33.340 393.355 34.700 ;
        RECT 4.000 27.180 393.755 33.340 ;
        RECT 4.400 25.820 393.755 27.180 ;
        RECT 4.400 25.180 393.355 25.820 ;
        RECT 4.000 23.820 393.355 25.180 ;
        RECT 4.000 19.020 393.755 23.820 ;
        RECT 4.400 17.020 393.755 19.020 ;
        RECT 4.000 16.300 393.755 17.020 ;
        RECT 4.000 14.300 393.355 16.300 ;
        RECT 4.000 9.500 393.755 14.300 ;
        RECT 4.400 8.140 393.755 9.500 ;
        RECT 4.400 7.500 393.355 8.140 ;
        RECT 4.000 6.975 393.355 7.500 ;
      LAYER met4 ;
        RECT 26.055 19.895 97.440 392.865 ;
        RECT 99.840 19.895 174.240 392.865 ;
        RECT 176.640 19.895 249.945 392.865 ;
  END
END wrapped_spraid
END LIBRARY

