VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_spraid
  CLASS BLOCK ;
  FOREIGN wrapped_spraid ;
  ORIGIN 0.000 0.000 ;
  SIZE 399.130 BY 409.850 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 405.850 53.870 409.850 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 69.100 399.130 70.300 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 0.000 257.190 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 0.000 269.150 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 0.000 79.630 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.390 0.000 397.950 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.430 0.000 385.990 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 0.000 128.390 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.820 4.000 73.020 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 168.380 399.130 169.580 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 105.820 399.130 107.020 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 0.000 281.110 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.790 405.850 163.350 409.850 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.150 0.000 354.710 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 277.180 399.130 278.380 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.070 405.850 102.630 409.850 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.790 405.850 347.350 409.850 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.300 4.000 335.500 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.630 405.850 372.190 409.850 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 405.850 218.550 409.850 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.070 0.000 263.630 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.270 0.000 226.830 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 405.850 121.030 409.850 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.270 405.850 65.830 409.850 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 405.850 144.950 409.850 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.590 0.000 361.150 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.030 0.000 183.590 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 86.780 399.130 87.980 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.030 405.850 22.590 409.850 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 249.980 399.130 251.180 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.430 0.000 293.990 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.860 4.000 398.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 0.000 116.430 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.670 0.000 153.230 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.990 0.000 287.550 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.020 4.000 100.220 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.620 4.000 45.820 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.550 405.850 304.110 409.850 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.390 0.000 305.950 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.430 405.850 316.990 409.850 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 213.260 399.130 214.460 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 313.900 399.130 315.100 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 205.100 399.130 206.300 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.580 4.000 162.780 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.070 0.000 171.630 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 405.850 365.750 409.850 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.500 4.000 90.700 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.030 0.000 367.590 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.900 4.000 9.100 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 0.000 98.030 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 368.300 399.130 369.500 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.830 405.850 335.390 409.850 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 0.000 30.870 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 0.000 109.990 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 195.580 399.130 196.780 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.830 0.000 220.390 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.420 4.000 154.620 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 405.850 213.030 409.850 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.500 4.000 362.700 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 405.850 84.230 409.850 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.030 405.850 390.590 409.850 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.270 405.850 249.830 409.850 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 341.100 399.130 342.300 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 349.260 399.130 350.460 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.180 4.000 244.380 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.350 405.850 340.910 409.850 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 232.300 399.130 233.500 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.030 405.850 114.590 409.850 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 59.580 399.130 60.780 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.380 4.000 407.580 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 405.850 90.670 409.850 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 376.460 399.130 377.660 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 160.220 399.130 161.420 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.460 4.000 207.660 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 405.850 35.470 409.850 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.420 4.000 18.620 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 0.000 190.030 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.750 405.850 267.310 409.850 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.550 405.850 396.110 409.850 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.780 4.000 325.980 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.830 0.000 36.390 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 405.850 181.750 409.850 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 32.380 399.130 33.580 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 405.850 353.790 409.850 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.580 4.000 26.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.620 4.000 181.820 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.950 0.000 299.510 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.590 405.850 384.150 409.850 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 405.850 285.710 409.850 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 222.780 399.130 223.980 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.660 4.000 370.860 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.190 0.000 342.750 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 133.020 399.130 134.220 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.230 405.850 261.790 409.850 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 405.850 310.550 409.850 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 78.620 399.130 79.820 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.100 4.000 36.300 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.630 405.850 280.190 409.850 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 405.850 139.430 409.850 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.070 405.850 194.630 409.850 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.830 405.850 243.390 409.850 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 0.000 336.310 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.180 4.000 108.380 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.550 0.000 373.110 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.230 0.000 54.790 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.380 4.000 271.580 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.390 405.850 236.950 409.850 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 141.180 399.130 142.380 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 14.700 399.130 15.900 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 405.850 40.990 409.850 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 331.580 399.130 332.780 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 397.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 397.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 397.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 397.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 397.360 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 405.850 169.790 409.850 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 395.500 399.130 396.700 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.980 4.000 353.180 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 240.460 399.130 241.660 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 322.060 399.130 323.260 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.060 4.000 289.260 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.430 0.000 17.990 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.270 0.000 134.830 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 41.900 399.130 43.100 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.870 405.850 231.430 409.850 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 0.000 158.750 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 6.540 399.130 7.740 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.230 0.000 330.790 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.510 405.850 17.070 409.850 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.260 4.000 316.460 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 187.420 399.130 188.620 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.700 4.000 389.900 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.100 4.000 172.300 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.350 0.000 317.910 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 405.850 157.830 409.850 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 0.000 140.350 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.660 4.000 234.860 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.100 4.000 308.300 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.900 4.000 145.100 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 405.850 151.390 409.850 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 0.000 104.470 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 405.850 96.190 409.850 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.990 0.000 379.550 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.870 0.000 208.430 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 304.380 399.130 305.580 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.780 4.000 53.980 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 0.000 86.070 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.910 405.850 127.470 409.850 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.030 0.000 275.590 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.580 4.000 298.780 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.390 405.850 328.950 409.850 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.830 405.850 59.390 409.850 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 405.850 132.990 409.850 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.630 405.850 188.190 409.850 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.670 405.850 176.230 409.850 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.910 0.000 12.470 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 0.000 61.230 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.380 4.000 135.580 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 0.000 165.190 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 385.980 399.130 387.180 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 405.850 72.270 409.850 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 405.850 224.990 409.850 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 0.000 42.830 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 96.300 399.130 97.500 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 286.700 399.130 287.900 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.500 4.000 226.700 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 177.900 399.130 179.100 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.070 405.850 10.630 409.850 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.980 4.000 81.180 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 358.780 399.130 359.980 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.790 405.850 255.350 409.850 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 0.000 91.590 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 113.980 399.130 115.180 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 0.000 245.230 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.950 0.000 391.510 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 405.850 29.030 409.850 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.830 0.000 312.390 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 0.000 49.270 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.230 0.000 146.790 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 51.420 399.130 52.620 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 403.660 399.130 404.860 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.220 4.000 127.420 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.790 0.000 324.350 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 123.500 399.130 124.700 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 0.000 6.030 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 294.860 399.130 296.060 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 405.850 377.710 409.850 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.630 0.000 349.190 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.750 405.850 359.310 409.850 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.860 4.000 262.060 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.900 4.000 281.100 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.390 0.000 213.950 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 0.000 250.750 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.460 4.000 343.660 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 405.850 77.790 409.850 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 405.850 206.590 409.850 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.700 4.000 253.900 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 0.000 67.670 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.870 0.000 24.430 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.190 405.850 273.750 409.850 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 405.850 200.150 409.850 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 0.000 177.150 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.950 405.850 322.510 409.850 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 24.220 399.130 25.420 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.180 4.000 380.380 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 267.660 399.130 268.860 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.630 0.000 73.190 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 0.000 122.870 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 0.000 195.550 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 259.500 399.130 260.700 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.430 0.000 201.990 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 405.850 298.590 409.850 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.590 405.850 292.150 409.850 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 405.850 47.430 409.850 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.510 405.850 109.070 409.850 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.230 0.000 238.790 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.630 405.850 4.190 409.850 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 395.130 150.700 399.130 151.900 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 397.295 404.175 ;
      LAYER met1 ;
        RECT 0.070 8.880 397.355 404.220 ;
      LAYER met2 ;
        RECT 0.100 405.570 3.350 407.165 ;
        RECT 4.470 405.570 9.790 407.165 ;
        RECT 10.910 405.570 16.230 407.165 ;
        RECT 17.350 405.570 21.750 407.165 ;
        RECT 22.870 405.570 28.190 407.165 ;
        RECT 29.310 405.570 34.630 407.165 ;
        RECT 35.750 405.570 40.150 407.165 ;
        RECT 41.270 405.570 46.590 407.165 ;
        RECT 47.710 405.570 53.030 407.165 ;
        RECT 54.150 405.570 58.550 407.165 ;
        RECT 59.670 405.570 64.990 407.165 ;
        RECT 66.110 405.570 71.430 407.165 ;
        RECT 72.550 405.570 76.950 407.165 ;
        RECT 78.070 405.570 83.390 407.165 ;
        RECT 84.510 405.570 89.830 407.165 ;
        RECT 90.950 405.570 95.350 407.165 ;
        RECT 96.470 405.570 101.790 407.165 ;
        RECT 102.910 405.570 108.230 407.165 ;
        RECT 109.350 405.570 113.750 407.165 ;
        RECT 114.870 405.570 120.190 407.165 ;
        RECT 121.310 405.570 126.630 407.165 ;
        RECT 127.750 405.570 132.150 407.165 ;
        RECT 133.270 405.570 138.590 407.165 ;
        RECT 139.710 405.570 144.110 407.165 ;
        RECT 145.230 405.570 150.550 407.165 ;
        RECT 151.670 405.570 156.990 407.165 ;
        RECT 158.110 405.570 162.510 407.165 ;
        RECT 163.630 405.570 168.950 407.165 ;
        RECT 170.070 405.570 175.390 407.165 ;
        RECT 176.510 405.570 180.910 407.165 ;
        RECT 182.030 405.570 187.350 407.165 ;
        RECT 188.470 405.570 193.790 407.165 ;
        RECT 194.910 405.570 199.310 407.165 ;
        RECT 200.430 405.570 205.750 407.165 ;
        RECT 206.870 405.570 212.190 407.165 ;
        RECT 213.310 405.570 217.710 407.165 ;
        RECT 218.830 405.570 224.150 407.165 ;
        RECT 225.270 405.570 230.590 407.165 ;
        RECT 231.710 405.570 236.110 407.165 ;
        RECT 237.230 405.570 242.550 407.165 ;
        RECT 243.670 405.570 248.990 407.165 ;
        RECT 250.110 405.570 254.510 407.165 ;
        RECT 255.630 405.570 260.950 407.165 ;
        RECT 262.070 405.570 266.470 407.165 ;
        RECT 267.590 405.570 272.910 407.165 ;
        RECT 274.030 405.570 279.350 407.165 ;
        RECT 280.470 405.570 284.870 407.165 ;
        RECT 285.990 405.570 291.310 407.165 ;
        RECT 292.430 405.570 297.750 407.165 ;
        RECT 298.870 405.570 303.270 407.165 ;
        RECT 304.390 405.570 309.710 407.165 ;
        RECT 310.830 405.570 316.150 407.165 ;
        RECT 317.270 405.570 321.670 407.165 ;
        RECT 322.790 405.570 328.110 407.165 ;
        RECT 329.230 405.570 334.550 407.165 ;
        RECT 335.670 405.570 340.070 407.165 ;
        RECT 341.190 405.570 346.510 407.165 ;
        RECT 347.630 405.570 352.950 407.165 ;
        RECT 354.070 405.570 358.470 407.165 ;
        RECT 359.590 405.570 364.910 407.165 ;
        RECT 366.030 405.570 371.350 407.165 ;
        RECT 372.470 405.570 376.870 407.165 ;
        RECT 377.990 405.570 383.310 407.165 ;
        RECT 384.430 405.570 389.750 407.165 ;
        RECT 390.870 405.570 395.270 407.165 ;
        RECT 0.100 4.280 395.960 405.570 ;
        RECT 0.790 4.000 5.190 4.280 ;
        RECT 6.310 4.000 11.630 4.280 ;
        RECT 12.750 4.000 17.150 4.280 ;
        RECT 18.270 4.000 23.590 4.280 ;
        RECT 24.710 4.000 30.030 4.280 ;
        RECT 31.150 4.000 35.550 4.280 ;
        RECT 36.670 4.000 41.990 4.280 ;
        RECT 43.110 4.000 48.430 4.280 ;
        RECT 49.550 4.000 53.950 4.280 ;
        RECT 55.070 4.000 60.390 4.280 ;
        RECT 61.510 4.000 66.830 4.280 ;
        RECT 67.950 4.000 72.350 4.280 ;
        RECT 73.470 4.000 78.790 4.280 ;
        RECT 79.910 4.000 85.230 4.280 ;
        RECT 86.350 4.000 90.750 4.280 ;
        RECT 91.870 4.000 97.190 4.280 ;
        RECT 98.310 4.000 103.630 4.280 ;
        RECT 104.750 4.000 109.150 4.280 ;
        RECT 110.270 4.000 115.590 4.280 ;
        RECT 116.710 4.000 122.030 4.280 ;
        RECT 123.150 4.000 127.550 4.280 ;
        RECT 128.670 4.000 133.990 4.280 ;
        RECT 135.110 4.000 139.510 4.280 ;
        RECT 140.630 4.000 145.950 4.280 ;
        RECT 147.070 4.000 152.390 4.280 ;
        RECT 153.510 4.000 157.910 4.280 ;
        RECT 159.030 4.000 164.350 4.280 ;
        RECT 165.470 4.000 170.790 4.280 ;
        RECT 171.910 4.000 176.310 4.280 ;
        RECT 177.430 4.000 182.750 4.280 ;
        RECT 183.870 4.000 189.190 4.280 ;
        RECT 190.310 4.000 194.710 4.280 ;
        RECT 195.830 4.000 201.150 4.280 ;
        RECT 202.270 4.000 207.590 4.280 ;
        RECT 208.710 4.000 213.110 4.280 ;
        RECT 214.230 4.000 219.550 4.280 ;
        RECT 220.670 4.000 225.990 4.280 ;
        RECT 227.110 4.000 231.510 4.280 ;
        RECT 232.630 4.000 237.950 4.280 ;
        RECT 239.070 4.000 244.390 4.280 ;
        RECT 245.510 4.000 249.910 4.280 ;
        RECT 251.030 4.000 256.350 4.280 ;
        RECT 257.470 4.000 262.790 4.280 ;
        RECT 263.910 4.000 268.310 4.280 ;
        RECT 269.430 4.000 274.750 4.280 ;
        RECT 275.870 4.000 280.270 4.280 ;
        RECT 281.390 4.000 286.710 4.280 ;
        RECT 287.830 4.000 293.150 4.280 ;
        RECT 294.270 4.000 298.670 4.280 ;
        RECT 299.790 4.000 305.110 4.280 ;
        RECT 306.230 4.000 311.550 4.280 ;
        RECT 312.670 4.000 317.070 4.280 ;
        RECT 318.190 4.000 323.510 4.280 ;
        RECT 324.630 4.000 329.950 4.280 ;
        RECT 331.070 4.000 335.470 4.280 ;
        RECT 336.590 4.000 341.910 4.280 ;
        RECT 343.030 4.000 348.350 4.280 ;
        RECT 349.470 4.000 353.870 4.280 ;
        RECT 354.990 4.000 360.310 4.280 ;
        RECT 361.430 4.000 366.750 4.280 ;
        RECT 367.870 4.000 372.270 4.280 ;
        RECT 373.390 4.000 378.710 4.280 ;
        RECT 379.830 4.000 385.150 4.280 ;
        RECT 386.270 4.000 390.670 4.280 ;
        RECT 391.790 4.000 395.960 4.280 ;
      LAYER met3 ;
        RECT 4.400 405.980 395.130 407.145 ;
        RECT 4.000 405.260 395.130 405.980 ;
        RECT 4.000 403.260 394.730 405.260 ;
        RECT 4.000 398.460 395.130 403.260 ;
        RECT 4.400 397.100 395.130 398.460 ;
        RECT 4.400 396.460 394.730 397.100 ;
        RECT 4.000 395.100 394.730 396.460 ;
        RECT 4.000 390.300 395.130 395.100 ;
        RECT 4.400 388.300 395.130 390.300 ;
        RECT 4.000 387.580 395.130 388.300 ;
        RECT 4.000 385.580 394.730 387.580 ;
        RECT 4.000 380.780 395.130 385.580 ;
        RECT 4.400 378.780 395.130 380.780 ;
        RECT 4.000 378.060 395.130 378.780 ;
        RECT 4.000 376.060 394.730 378.060 ;
        RECT 4.000 371.260 395.130 376.060 ;
        RECT 4.400 369.900 395.130 371.260 ;
        RECT 4.400 369.260 394.730 369.900 ;
        RECT 4.000 367.900 394.730 369.260 ;
        RECT 4.000 363.100 395.130 367.900 ;
        RECT 4.400 361.100 395.130 363.100 ;
        RECT 4.000 360.380 395.130 361.100 ;
        RECT 4.000 358.380 394.730 360.380 ;
        RECT 4.000 353.580 395.130 358.380 ;
        RECT 4.400 351.580 395.130 353.580 ;
        RECT 4.000 350.860 395.130 351.580 ;
        RECT 4.000 348.860 394.730 350.860 ;
        RECT 4.000 344.060 395.130 348.860 ;
        RECT 4.400 342.700 395.130 344.060 ;
        RECT 4.400 342.060 394.730 342.700 ;
        RECT 4.000 340.700 394.730 342.060 ;
        RECT 4.000 335.900 395.130 340.700 ;
        RECT 4.400 333.900 395.130 335.900 ;
        RECT 4.000 333.180 395.130 333.900 ;
        RECT 4.000 331.180 394.730 333.180 ;
        RECT 4.000 326.380 395.130 331.180 ;
        RECT 4.400 324.380 395.130 326.380 ;
        RECT 4.000 323.660 395.130 324.380 ;
        RECT 4.000 321.660 394.730 323.660 ;
        RECT 4.000 316.860 395.130 321.660 ;
        RECT 4.400 315.500 395.130 316.860 ;
        RECT 4.400 314.860 394.730 315.500 ;
        RECT 4.000 313.500 394.730 314.860 ;
        RECT 4.000 308.700 395.130 313.500 ;
        RECT 4.400 306.700 395.130 308.700 ;
        RECT 4.000 305.980 395.130 306.700 ;
        RECT 4.000 303.980 394.730 305.980 ;
        RECT 4.000 299.180 395.130 303.980 ;
        RECT 4.400 297.180 395.130 299.180 ;
        RECT 4.000 296.460 395.130 297.180 ;
        RECT 4.000 294.460 394.730 296.460 ;
        RECT 4.000 289.660 395.130 294.460 ;
        RECT 4.400 288.300 395.130 289.660 ;
        RECT 4.400 287.660 394.730 288.300 ;
        RECT 4.000 286.300 394.730 287.660 ;
        RECT 4.000 281.500 395.130 286.300 ;
        RECT 4.400 279.500 395.130 281.500 ;
        RECT 4.000 278.780 395.130 279.500 ;
        RECT 4.000 276.780 394.730 278.780 ;
        RECT 4.000 271.980 395.130 276.780 ;
        RECT 4.400 269.980 395.130 271.980 ;
        RECT 4.000 269.260 395.130 269.980 ;
        RECT 4.000 267.260 394.730 269.260 ;
        RECT 4.000 262.460 395.130 267.260 ;
        RECT 4.400 261.100 395.130 262.460 ;
        RECT 4.400 260.460 394.730 261.100 ;
        RECT 4.000 259.100 394.730 260.460 ;
        RECT 4.000 254.300 395.130 259.100 ;
        RECT 4.400 252.300 395.130 254.300 ;
        RECT 4.000 251.580 395.130 252.300 ;
        RECT 4.000 249.580 394.730 251.580 ;
        RECT 4.000 244.780 395.130 249.580 ;
        RECT 4.400 242.780 395.130 244.780 ;
        RECT 4.000 242.060 395.130 242.780 ;
        RECT 4.000 240.060 394.730 242.060 ;
        RECT 4.000 235.260 395.130 240.060 ;
        RECT 4.400 233.900 395.130 235.260 ;
        RECT 4.400 233.260 394.730 233.900 ;
        RECT 4.000 231.900 394.730 233.260 ;
        RECT 4.000 227.100 395.130 231.900 ;
        RECT 4.400 225.100 395.130 227.100 ;
        RECT 4.000 224.380 395.130 225.100 ;
        RECT 4.000 222.380 394.730 224.380 ;
        RECT 4.000 217.580 395.130 222.380 ;
        RECT 4.400 215.580 395.130 217.580 ;
        RECT 4.000 214.860 395.130 215.580 ;
        RECT 4.000 212.860 394.730 214.860 ;
        RECT 4.000 208.060 395.130 212.860 ;
        RECT 4.400 206.700 395.130 208.060 ;
        RECT 4.400 206.060 394.730 206.700 ;
        RECT 4.000 204.700 394.730 206.060 ;
        RECT 4.000 199.900 395.130 204.700 ;
        RECT 4.400 197.900 395.130 199.900 ;
        RECT 4.000 197.180 395.130 197.900 ;
        RECT 4.000 195.180 394.730 197.180 ;
        RECT 4.000 190.380 395.130 195.180 ;
        RECT 4.400 189.020 395.130 190.380 ;
        RECT 4.400 188.380 394.730 189.020 ;
        RECT 4.000 187.020 394.730 188.380 ;
        RECT 4.000 182.220 395.130 187.020 ;
        RECT 4.400 180.220 395.130 182.220 ;
        RECT 4.000 179.500 395.130 180.220 ;
        RECT 4.000 177.500 394.730 179.500 ;
        RECT 4.000 172.700 395.130 177.500 ;
        RECT 4.400 170.700 395.130 172.700 ;
        RECT 4.000 169.980 395.130 170.700 ;
        RECT 4.000 167.980 394.730 169.980 ;
        RECT 4.000 163.180 395.130 167.980 ;
        RECT 4.400 161.820 395.130 163.180 ;
        RECT 4.400 161.180 394.730 161.820 ;
        RECT 4.000 159.820 394.730 161.180 ;
        RECT 4.000 155.020 395.130 159.820 ;
        RECT 4.400 153.020 395.130 155.020 ;
        RECT 4.000 152.300 395.130 153.020 ;
        RECT 4.000 150.300 394.730 152.300 ;
        RECT 4.000 145.500 395.130 150.300 ;
        RECT 4.400 143.500 395.130 145.500 ;
        RECT 4.000 142.780 395.130 143.500 ;
        RECT 4.000 140.780 394.730 142.780 ;
        RECT 4.000 135.980 395.130 140.780 ;
        RECT 4.400 134.620 395.130 135.980 ;
        RECT 4.400 133.980 394.730 134.620 ;
        RECT 4.000 132.620 394.730 133.980 ;
        RECT 4.000 127.820 395.130 132.620 ;
        RECT 4.400 125.820 395.130 127.820 ;
        RECT 4.000 125.100 395.130 125.820 ;
        RECT 4.000 123.100 394.730 125.100 ;
        RECT 4.000 118.300 395.130 123.100 ;
        RECT 4.400 116.300 395.130 118.300 ;
        RECT 4.000 115.580 395.130 116.300 ;
        RECT 4.000 113.580 394.730 115.580 ;
        RECT 4.000 108.780 395.130 113.580 ;
        RECT 4.400 107.420 395.130 108.780 ;
        RECT 4.400 106.780 394.730 107.420 ;
        RECT 4.000 105.420 394.730 106.780 ;
        RECT 4.000 100.620 395.130 105.420 ;
        RECT 4.400 98.620 395.130 100.620 ;
        RECT 4.000 97.900 395.130 98.620 ;
        RECT 4.000 95.900 394.730 97.900 ;
        RECT 4.000 91.100 395.130 95.900 ;
        RECT 4.400 89.100 395.130 91.100 ;
        RECT 4.000 88.380 395.130 89.100 ;
        RECT 4.000 86.380 394.730 88.380 ;
        RECT 4.000 81.580 395.130 86.380 ;
        RECT 4.400 80.220 395.130 81.580 ;
        RECT 4.400 79.580 394.730 80.220 ;
        RECT 4.000 78.220 394.730 79.580 ;
        RECT 4.000 73.420 395.130 78.220 ;
        RECT 4.400 71.420 395.130 73.420 ;
        RECT 4.000 70.700 395.130 71.420 ;
        RECT 4.000 68.700 394.730 70.700 ;
        RECT 4.000 63.900 395.130 68.700 ;
        RECT 4.400 61.900 395.130 63.900 ;
        RECT 4.000 61.180 395.130 61.900 ;
        RECT 4.000 59.180 394.730 61.180 ;
        RECT 4.000 54.380 395.130 59.180 ;
        RECT 4.400 53.020 395.130 54.380 ;
        RECT 4.400 52.380 394.730 53.020 ;
        RECT 4.000 51.020 394.730 52.380 ;
        RECT 4.000 46.220 395.130 51.020 ;
        RECT 4.400 44.220 395.130 46.220 ;
        RECT 4.000 43.500 395.130 44.220 ;
        RECT 4.000 41.500 394.730 43.500 ;
        RECT 4.000 36.700 395.130 41.500 ;
        RECT 4.400 34.700 395.130 36.700 ;
        RECT 4.000 33.980 395.130 34.700 ;
        RECT 4.000 31.980 394.730 33.980 ;
        RECT 4.000 27.180 395.130 31.980 ;
        RECT 4.400 25.820 395.130 27.180 ;
        RECT 4.400 25.180 394.730 25.820 ;
        RECT 4.000 23.820 394.730 25.180 ;
        RECT 4.000 19.020 395.130 23.820 ;
        RECT 4.400 17.020 395.130 19.020 ;
        RECT 4.000 16.300 395.130 17.020 ;
        RECT 4.000 14.300 394.730 16.300 ;
        RECT 4.000 9.500 395.130 14.300 ;
        RECT 4.400 8.140 395.130 9.500 ;
        RECT 4.400 7.500 394.730 8.140 ;
        RECT 4.000 6.975 394.730 7.500 ;
      LAYER met4 ;
        RECT 96.895 11.735 97.440 286.785 ;
        RECT 99.840 11.735 174.240 286.785 ;
        RECT 176.640 11.735 251.040 286.785 ;
        RECT 253.440 11.735 327.840 286.785 ;
        RECT 330.240 11.735 343.785 286.785 ;
  END
END wrapped_spraid
END LIBRARY

